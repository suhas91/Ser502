var stackVar = STACK;

print "push element onto stack";
stackVar.push(1);

print "push element onto stack";
stackVar.push(2);

print "push element onto stack";
stackVar.push(3);

print "push element onto stack";
stackVar.push(4);

print "push element onto stack";
stackVar.push(5);

print "push element onto stack";
stackVar.push(6);

print "push element onto stack";
stackVar.push(7);

print "push element onto stack";
stackVar.push(8);

print "push element onto stack";
stackVar.push(9);

print "push element onto stack";
stackVar.push(10);

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;

print "element popped";
popEle = stackVar.pop();
print popEle;