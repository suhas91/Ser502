var x = 5;
var y = 10;

if( x == y ){
	print "entered if block";
	print x;
	print "both are equal";
} else{
	print "both the numers are unequal";
}