 var num = 10;
 
while( num > 1 ){
	print num;
	num = num-1;
}
print "exited while loop";